00a29403
403402b3
001404b3
